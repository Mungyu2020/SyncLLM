

module Q3bFSM
(
  input clk,
  input reset,
  input x,
  output z
);

  parameter A = 0;parameter B = 1;parameter C = 2;parameter D = 3;parameter E = 4;
  reg [2:0] state;reg [2:0] next_state;

  always @(posedge clk) begin
    if(reset) state <= A; 
    else state <= next_state;
  end


  always @(*) begin
    case(state)
      A: next_state <= (x)? B : A;
      B: next_state <= (x)? E : B;
      C: next_state <= (x)? B : C;
      D: next_state <= (x)? C : B;
      E: next_state <= (x)? E : D;
      default: next_state <= A;
    endcase
  end

  assign z = (state == D) || (state == E);

endmodule

